--ola